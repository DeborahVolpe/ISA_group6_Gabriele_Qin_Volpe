library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;

entity data_sink is
  port (
    CLK   : in std_logic;  -- clock signal
    RST_n : in std_logic; --reset low active
    VIN   : in std_logic; -- valid output of the filter
    DIN   : in signed(10 downto 0) -- output of the IIR filter
	);
end data_sink;

architecture beh of data_sink is

begin  -- beh

  process (CLK, RST_n)
    file res_fp : text open WRITE_MODE is "./results.txt";
    variable line_out : line;    
  begin  -- process
    if RST_n = '0' then                 -- asynchronous reset (active low)
      null;
    elsif CLK'event and CLK = '1' then  -- rising clock edge
      if (VIN = '1') then
        write(line_out, to_integer(DIN));
        writeline(res_fp, line_out);
      end if;
    end if;
  end process;

end beh;
